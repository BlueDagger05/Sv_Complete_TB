package apb_states;
	typedef enum logic [1:0] {IDLE, SETUP, ACCESS} apb_states;
endpackage: apb_states
