package checker_pkg;
	import apb_slave_ifc::*;
	
class Checker;
	
	
endclass: Checker	
endpackage : checker_pkg